/*
Digital thermometer reads off temperature from temperature sensor with I2C interface
and sends data to PC over UART. PC displays data on console.

Additionally PC can send write/read requests to temperature sensor.
Options include reading 1/2 bytes or writing 1 or 2 bytes to 
temperature registers/status registers or configuration registers.

Since all functionality of temperature sensor is implemented in terms of reads/writes to its
registers further info can be found on the temperature sensor's datasheet (ADT7420)

On PC side, user types in the instruction and the corresponding data is sent to the FPGA 
through UART. Transmission requires that the data comes in the packet : 
-Start Byte: 8 bit signal all bits high to indicate start of instruction
-Address Byte: address of register on temperature sensor to which operation is directed
-Operation Byte: operation to be performed (read/write)
-(Optional) Data Byte 1: Byte/LSB to be written to temperature register
-(Optional) Data Byte 2: Byte/MSB to be written to temperature register
-Stop Byte: 8-bit signal all bits high to indicate end of instruction.

Should the user delay in sending the necessary instruction in full, then
a grace period of 10 seconds is given before a the system times out and the
user is required to retype the instruction in its entirety.

Buffers are added to store the instruction's as they await execution by the
I2C controller. Buffers are also added to store the results of the I2C transaction.

If buffers fill up, 8 led's light up indicating that the buffers are full.
Hence users should retype their instructions when buffers are full and
refrain from sending in too many instructions at once.

*/



module temp_sensor (input logic clk,reset,
				   	input logic tx, //Data bit from PC UART transmitter
				    input logic sample_tick, //Sample_tick from baud rate generator
				    input logic[9:0] dvsr, //Adjust UART and I2C frequency using FPGA slide switches
				    output logic[7:0] data_byte, //Data byte transmitted to UART.
				    output logic[15:0] led_on,
				    output tri scl, //SCL is I2C clock generated by I2C controller and SDA is I2C data line
				    inout tri sda);
				    
				    logic time_out, buffers_full ;//If there is more than 10 seconds delay in typing in instructions or in case too many instructions are being sent.
				    	    
				    	    
				    	    
				    logic rx_done_tick;
				    logic[7:0] received_byte_next,received_byte_reg;
				    	   
				    	    
				    uart_rx uart_receiver(.*,
				    	    			  .rx_done_tick(rx_done_tick),
				    	    			  .received_byte(received_byte_next));
				    	    
				    	    logic valid;
				    	    logic rx_done;
				    	    
				    	    logic waiting;
				    	    
				    	    //TIME_OUT AND TEMP SENSOR BUSY LED REGISTER
				    	    always_ff @(posedge clk, posedge reset) 
				    	    	if(reset) begin
				    	    		led_on <= '0;
				    	    	end
				    	    	
				    	    	else begin
				    	    		led_on[0] <= waiting;
				    	    		led_on[7:1] <= (time_out) ? '1:'0;
				    	    		led_on[15:8] <= (buffers_full) ? '1:'0;
				    	    	end
				    	    	
				    	    //UART - UART-I2C BRIDGE INTERFACE REGISTER
				    	    always_ff @(posedge clk, posedge reset)
				    	    	if(reset) begin
				    	    		rx_done <= '0;
				    	    		received_byte_reg <= '0;
				    	    	end
				    	    	
				    	    	else begin
				    	    		rx_done <= rx_done_tick;
				    	    		received_byte_reg <= received_byte_next;
				    	    	end
				    	
				    	     /*Indicates availability of I2C controller for initiating another I2C transaction. 
				    	     Controller becomes available as soon as it sends off acquired data to I2C-UART stage provided
				    	     I2C-UART stage isn't stacked with previous requests awaiting transmission.
				    	     */
				    	     logic initiate, initiate_next;
				    	     logic i2c_ready; 
				    	     logic[2:0] mode, mode_next;
				    	     logic[7:0] addr_pointer, addr_pointer_next;
				    	     logic[15:0] wr_data, wr_data_next;
				    	     
				    	     logic wr_databuffer1, wr_databuffer2, wr_opbuffer,wr_addrbuffer;
				    	     logic wr_databuffer1_next, wr_databuffer2_next, wr_opbuffer_next,wr_addrbuffer_next;
				    	   
				    	   //All 3 signals above are commands and data sent to i2c core.
				    	     uart_i2c_tramsmitter uart_i2c_bridge(.*,
				    	     										.time_out(time_out),
				    	     										.buffers_full(buffers_full),
				    	     										.waiting(waiting),
				    	    										.initiate(initiate_next),
				    	    										.received_byte(received_byte),
				    	    										.rx_done_tick(rx_done),
				    	    										.i2c_ready(i2c_ready),
				    	    										.mode(mode_next),
				    	    										.addr_pointer(addr_pointer_next),
				    	    										.wr_data(wr_data_next),
				    	    										.wr_addrbuffer(wr_addrbuffer_next),
				    	    										.wr_databuffer1(wr_databuffer1_next),
				    	    										.wr_databuffer2(wr_databuffer2_next),
				    	    										.wr_opbuffer(wr_opbuffer_next));
				    	    	
				    	    	
				    	    	//UART-I2C TRANSMITTER TO I2C WAIT STAGE REGISTER
				    	    	always_ff @(posedge clk,posedge reset)
				    	    		if(reset) begin
				    	    			wr_addrbuffer <= '0;
				    	    			wr_databuffer1 <= '0;
				    	    			wr_databuffer2 <= '0;
				    	                        wr_opbuffer <= '0;
				    	                        addr_pointer <= '0;
				    	                        mode <= '0;
				    	                        wr_data <= '0;
				    	                        initiate <= '0;
				    	                end
				    	                
				    	                else begin
				    	                	wr_addrbuffer <= wr_addrbuffer_next;
				    	                	wr_databuffer1 <= wr_databuffer1_next;
				    	                	wr_databuffer2 <= wr_databuffer2_next;
				    	                	wr_opbuffer <= wr_opbuffer_next;
				    	                	addr_pointer <= addr_pointer_next;
				    	                	wr_data <= wr_data_next;
				    	                	mode <= mode_next;
				    	                	initiate <= initiate_next;
				    	                end
				    	                
				    	                
				    	        //Logic to determine what data is passed to I2C controller
				    	    	//Signals on output of register remain the same unless we initiate a new write if not we initiate continous read operation.
				    	    	logic[15:0] i2c_data;
				    	    	logic[7:0] i2c_address;
				    	    	logic[2:0] i2c_op;
				    	    	logic[1:0] valid_instr; //Use lower bit as an initiate signal for i2c transaction and upper bit as indication of whether instruction is non-queried(0 for non-queried)
				    	    	logic transmit_complete; //Has I2C data been transmitted to PC.
				    	                
				    	        uart_i2c_arbiter uart_to_i2c(.*,
				    	        							.i2c_data(i2c_data),
				    	        							.i2c_op(i2c_op),
				    	        							.valid_instr(valid_instr),
				    	        							.i2c_address(i2c_address),
				    	        							.transmit_complete(transmit_complete),
				    	        							.i2c_ready(i2c_ready),
				    	        							.initiate(initiate),
				    	        							.wr_addrbuffer(wr_addrbuffer),
				    	        							.wr_databuffer1(wr_databuffer1),
				    	        							.wr_databuffer2(wr_databuffer2),
				    	        							.wr_opbuffer(wr_opbuffer),
				    	        							.addr_pointer(addr_pointer),
				    	        							.wr_data(wr_data),
				    	        							.mode(mode));
				    	        
				    	        
				    	                        
				    	    			
				    	    			
				    	    	logic[15:0] i2c_rx_data_next, i2c_rx_data_reg;
				    	    	logic i2c_data_rdy, i2c_data_rdy_next;
				    	    	logic[3:0] fail_signals_next, fail_signals_reg;
				    	    	logic default_mode_next, default_mode_reg;
				    	    	logic i2c_ready_reg, i2c_ready_next;
				    	    	logic full_i2c_databuffer;
				    	    	i2cmaster i2ccontroller(.*,
				    	    						       .full_i2cdatabuffer(full_i2cdatabuffer),
				    	    						       .wr_data(i2c_data),
				    	    						       .initiate(valid_instr[0]),
				    	    						       .is_default_op(valid_instr[1]),
				    	    						       .mode(i2c_op),
				    	    						       .serialbusaddr(7'b1001000),
				    	    						       .addrpointer(i2c_address),
				    	    						       .received_data(i2c_rx_data_next),
				    	    						       .ready(i2c_ready_next),
				    	    						       .continous_mode_output(default_mode_next),
				    	    						       .i2c_data_rdy(i2c_data_rdy_next),
				    	    						       .failure_signal(fail_signals_next));
				    	    	
				    	    	
				    	    	//Register in between I2C controller and I2C - UART ARBITER STAGE
				    	    	always_ff @(posedge clk, posedge reset) 
				    	    		if(reset) begin
				    	    			i2c_rx_data_reg <= '0;
				    	    			fail_signals_reg <= '0;
				    	    			default_mode_reg <= '0;
				    	    			i2c_ready_reg <= '0;
				    	    			i2c_data_rdy <= '0;
				    	    		end
				    	    		
				    	    		else begin
				    	    			i2c_rx_data_reg <= i2c_rx_data_next;
				    	    			fail_signals_reg <= fail_signals_next;
				    	    			default_mode_reg <= default_mode_next;
				    	    			i2c_ready_reg <= i2c_ready_next;
				    	    			i2c_data_rdy <= i2c_data_rdy_next;
				    	    		end
				    	    		
				    	    		
				    	    	
				    	    	//I2C-uart arbitrer. Determine whether UART transmission can take place depending on data info. Results asked for take priority.
				    	    			
				    	    			
				
				     	logic[15:0] toPC_data;
				     	logic[7:0] toPC_address;
				     	logic[7:0] toPC_mode;
				     	logic data_rdy;
				     
				     	i2c_uart_arbiter i2c_to_uart (.*,
				     								 .toPC_data(toPC_data),
				     								 .toPC_address(toPC_address),
				     								 .toPC_mode(toPC_mode),
				     								 .data_ready(data_rdy), //Output signal that indicates whether data is ready for transmission
				     								 .i2c_rx_data(i2c_rx_data_reg),
				     								 .addr_pointer(addr_pointer_next),
				     								 .mode(mode_next),
				     								 .default_mode(default_mode_reg),
				     								 .i2c_data_rdy(i2c_data_rdy),
				     								 .transmit_complete(transmit_complete),
				     								 .fail_signals(fail_signals_reg),
				     								 .full_i2cdatabuffer(full_i2cdatabuffer));
				     	
				     	//i2c to uart arbiter has register for passing data to i2c-uart bridge built in. Thus we need only make direct connections
				     	
				    	
				    	logic[7:0] tx_byte, tx_byte_next;
				    	logic tx_start, tx_start_next; //Get UART to start transmission 
				    	logic tx_done_tick, tx_done_tick_next; //UART indication that it finished sending the byte
				    	
				    	//For your own sake have internal registers that store the necessary data bytes.
				        i2c_uart_transmitter i2c_uart_bridge (.*,
				    	    									  .data_ready(data_rdy),
				    	    									  .tx_done_tick(tx_done_tick),
				    	    									  .received_data(toPC_Data),
				    	    									  .op_data(toPC_mode),
				    	    									  .addr_pointer(toPC_address),
				    	    									  .tx_start(tx_start_next),
				    	    									  .data_byte(tx_byte_next),
				    	    									  .transmit_complete(transmit_complete));
				    	    									  
				    	
				    	//Intermediary register
				    	always_ff @(posedge clk, posedge reset)
				    		if(reset) begin
				    			tx_byte <= '0;
				    			tx_start <= '0;
				    			tx_done_tick <= '0;
				    		end
				    		
				    		else begin
				    			tx_byte <= tx_byte_next;
				    			tx_start <= tx_start_next;
				    			tx_done_tick <= tx_done_tick_next;
				    		end
				    		
				    	
				    	uart_tx uart_transmitter(.*,
				    							 .data_byte(tx_byte),
				    							 .tx_start(tx_start),
				    							 .tx_done_tick(tx_done_tick_next));
				    							 
				    	
endmodule  
