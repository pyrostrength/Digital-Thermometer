/*I2c controller works for reading and writing bytes to i2c temp sensor*/

module i2cmaster_test ;
    
    ////INPUTS
    logic clk,reset;
    
    /*If buffers on next pipeline stage are full,
    we do not initiate communication*/
	logic full_i2cbuffer; 
	//Data to write to temp sensor registers
	logic[15:0] wr_data;
	
	/*Operation to be performed. 1st 4 bits
	are {write_2byte, write_1byte,read_2byte,read_1byte}*/
	logic[7:0] mode;
	
	//signal to initiate I2C communication
	logic[1:0] valid_instr;
	
	//address of temperature sensor registe			 
	logic[7:0] reg_address;
	////INPUTS
	
	////OUTPUTS
	//Indicates controller is ready to initiate communication
	logic master_free; 
	
	//Indicates read/write failure
	logic[6:0] failure_signal;
	
	//Indicates completion of communication
	logic i2c_data_rdy;
				 
	/*Info for completed instruction to be passed onto next pipeline
	stage*/
	logic[1:0] i2c_valid_instr;
	
	logic[15:0] i2c_retrieved_data;
	
	logic[7:0] i2c_op_info;
	
	logic[7:0] i2c_instr_address;
				 
	wire scl; //SCL clock generated by master
	
	
	//Actual SDA line
	wire SDA; //Serial Data Line.
	////OUTPUTS
	
	
	logic[6:0] serialbusaddr;
	
	assign serialbusaddr = 7'b1001000;
	
	//Holds data byte to be written by I2C controller
	logic[8:0] write_vector;
	
	//Indicates failure to receive ack or nack bit
	logic send_fail;
	
	typedef enum { 
				    idle,start1,start2, address1,address2,address3,address4,address5,address6,
				    restart1,restart2,restart3,restart4,
				    read1,read2,read3,read4,read5,read6,
				    write1,write2,write3,write4,write5,write6,
				    stop1,stop2,stop3} state_type;
	
	i2cmaster #(.SYS_CLK_FREQ(100000000),.SCL_FREQ(3000000)) controller(.*,
	                                                                   .sda(SDA));
	
	/*Let sda_reg represent the value that slave 
	drives the wire sda. Wire sda is connected to
	tri-state buffer in controller*/
	logic sda_reg;
	
	/*SDA line has a pullup resistor connected to it
	thus it's driven high when output on master or 
	slave is in high impedance state*/
	/*sda_reg is driving signal of slave device*/
	assign (highz1,strong0) SDA = sda_reg;
	
	/*sda is driving signal for master device*/
	//assign (highz1,strong0) SDA = sda;
	
	/*model of pullup resistor on sda line*/
	assign (pull1,strong0) SDA = 1'b1;
	
	/*model of pullup resistor on scl line*/
	assign (pull1,strong0) scl = 1'b1;
	
	int dvsr = (100000000/3000000);
	/*Provides the number of system clock cycles per a third of SCL period. Although  
	integer division may round down or up we need not worry about this in
	simulation as design accounts for it*/
	int third = (100000000/(3000000*3)); 
	
	`timescale 1ns/1ps
	
	always begin
		#5 clk = ~clk;
	end
	
	
	/*Task randomizes the data inputs for 
	transmission.
	*/
	task automatic randomized_inputs;
	   output logic[1:0] valid;
	   output logic full_buffer;
	   output logic[15:0] data;
	   output logic[7:0] mode;
	   output logic[7:0] address;
	   
	   /*Create a logic vector that runs
	   from 0 to 3. Operation info encoded
	   in a 7 bit 1 hot signal*/
	   automatic logic[1:0] bit_pos;
	   
	   /*Randomize operation to be performed*/
	   bit_pos = $random();
	   
	   begin
	       /*Note that mode may be read but
	       data value returned is a non-zero
	       number. Thus we must ensure
	       that if mode is read/write byte we don't load*/
	       
	       full_buffer = $random();
	       valid = $random();
	       data = $random();
	       mode = 8'b0000_0001 << bit_pos;
	       address = $random();
	      
	   end
	endtask
	
	
	/*Tasks for checking that correct data bit is
	placed on sda line by controller when it writes
	bytes such as the serial bus address, register
	address or data bytes. Also checks to see if
	ack/nack bit is received and whether failure signal
	is asserted.
	
	Must pass data byte to be placed on sda and through int
	k indicate which failure signal to look at
	Recall failure signal vector format is
	{sba_send_fail, address_send_fail, write_byte1_fail, 
	write_byte2_fail, read_byte1_fail, read_byte2_fail}*/
	task automatic write_phase_check;
	   input logic[9:0] write_vector;
	   input int k;
	   logic val;
	   
	   //Bit to write on SDA
	   //logic write_bit;
	   //In last half of SCL low phase
	   for (int i = 0; i < 9; i++) begin
	       //sda_reg = (i == 8) ? 'z:'0;
	       //write_bit = (i<8) ? write_vector[8-i] : sda_reg;
	       
	       assert(scl == '0) begin
		   end else begin $display("SCL not pulled low before writing to SDA");
		   end
		      
		   //Write phase before receiving ack/nack bit
		   if(i < 8) begin
		      assert(SDA == write_vector[8-i]) begin
		      end else begin 
		      $display("Appropriate bit not shifted out");
		      $display("error is here");
		      $display(write_vector[8-i]);
		      $display(SDA);
		      end
		   end
		      
		   else begin
		      //Randomize the received ack bit
		      val = $random(); //Randomize the received ack bit
		      if (val == '0) begin
		      //Received the ack bit
		          sda_reg = val;
		          send_fail = '0;
		      end
		      
		      //Haven't received the appropriate ack bit
		      else if(val != '0) begin
		          sda_reg = 'z;
		          send_fail = '1;
		      end
		   end
		      
		   #((third)*10);
		      
		   /*High phase of SCL clock during which
		   sda line is sampled even when controller is
		   writing to sda line. Thus for each byte written
		   by the controller, the byte written is stored in
		   a register.*/
		      
		   assert(scl == '1) begin
		   end else begin 
		   $display("SCL clock not high");
		   $display($time);
		   end
		      
		   /*Output data bits during writes
		   is always the most significant bit of a vector
		   left shifted by 1 bit for every bit sent.
		   We sample data on SDA at the end of SCL high
		   phase so we shall make the check on the
		   subsequent low phase*/
		   if(i < 8) begin
		      assert(SDA == write_vector[8-i]) begin
		      end else begin 
		      $display("Appropriate bit not shifted out");
		      $display("error is here");
		      end
		   end
		   
		   /*Regardless sda line should be driven by slave*/
		   else begin
		      assert(SDA == val) begin
		      end else begin $display("SDA not driven by slave");
		      end
		   end
		      
		   #((third)*10);
		      
		   /*Low phase of SCL clock during which
		   we check for send failure. Recall that sda line is
		   driven by slave in the final loop iteration*/
		   assert(scl == '0) begin
		   end else begin 
		   $display("SCL clock not low prior to next data bit transfer");
		   $display($time);
		   
		   end
		      
		   if(i < 8) begin
		      assert(SDA == write_vector[8-i]) begin
		      end else begin 
		      $display("Appropriate bit not shifted out");
		      end
		   end
		   
		   else begin
		      /*Ensure operation success or failure was recorded*/
		      assert(failure_signal[k] == send_fail) begin
		      end else begin $display("Success or failure of operation not indicated properly");
		      end
		      
		      /*Ensure sda line is driven by slave */
		      assert(SDA == val) begin
		      end else begin $display("SDA not driven by slave");
		      end
		   end
		   
		   //Slave lets go of SDA during low phase
		   #((third-1)*10);
		   
		   sda_reg = 'z;
		   #10;  
		end    
	endtask
	
	/*For read operations, after sending register address
	byte a repeat start is initiated, then the serial bus
	address is sent + a high bit then the data bytes are
	read. If 1 byte is read a nack is sent from master. If
	2 bytes a read an ack is sent by master after the first byte 
	and a nack after the second byte. We then proceed to the stop
	state*/
	task automatic read_phase_check;
	   input logic[7:0] mode;
	   /*We randomize the data byte
	   that will be read from temp sensor*/
	   output logic [1:0][7:0] databyte;
	   int count,k;
	   databyte = $random();
	   
	   /*We run thru the loop twice if
	   reading 2 bytes but once if reading
	   1 byte*/
	   count = (mode[1]) ? 2:1;
	   /*We first initiate the repeat start*/
	   //In restart 1 state where SDA has been pulled high
	   assert(SDA == '1) begin
	   end else begin $display("SDA hasn't been pulled high before restart");
	   end
	   
	   assert(scl == '0) begin
	   end else begin $display("SCL should start low before restart");
	   end
	   
	   #(third*10);
	   
	   //In restart 2 state
	   assert(SDA == '1) begin
	   end else begin $display("SDA should be high as SCL high for restart");
	   end
	   
	   assert(scl == '1) begin
	   end else begin $display("SCL should be high");
	   end
	   
	   #(third*10);
	   
	   //In restart 3 state
	   assert(SDA == '0) begin
	   end else begin $display("SDA should be low to signal new start");
	   end
	   
	   assert(scl == '1) begin
	   end else begin $display("SCL should be high with SDA falling to signal new start");
	   end
	   
	   #(third*10);
	   //In restart 4 state
	   assert(SDA == '0) begin
	   end else begin $display("SDA should be low to finalize restart");
	   end 
	   
	   assert(scl == '0) begin
	   end else begin $display("scl should be low to finalize restart");
	   end
	   
	   #(third*10);
	   /*We then write serial bus address byte
	   and an active high signal to temp sensor*/
	   write_vector = {serialbusaddr, 1'b1, '0};
	   write_phase_check(write_vector,2);
	   
	   //Transition into read state 
	   /*Loop iterator variable*/
	   k = 0;
	   while(k < count) begin
	       /*Loop iterates thru all the bits
	       transmitted in a single frame*/
	       for(int i = 0; i<9 ; i++) begin
	           /*Reading the byte*/
	           if(i<8) begin
	               /*Most significant bit of
	               most significant byte is shifted out
	               first*/
	               sda_reg = databyte[1-k][7-i];
	               
	               #10;
	               
	               assert(SDA == sda_reg) begin
	               end else begin $display("Slave hasn't taken control of SDA line during read");
	               end
	               
	               assert(scl == '0) begin
	               end else begin $display("SCL line isn't low when new read data received");
	               end
	               
	               #((third-1)*10);
	               //Read 2 state
	               
	               assert(SDA == sda_reg) begin
	               end else begin 
	               $display("Slave has changed SDA control during SCL high phase");
	               end
	               
	               assert(scl == '1) begin
	               end else begin $display("SCL line isn't high");
	               end
	               
	               #(third*10);
	               //Read 3 state
	               assert(SDA == sda_reg) begin
	               end else begin 
	               $display("Slave has changed SDA control during SCL low phase");
	               end
	               
	               assert(scl == '0) begin
	               end else begin $display("SCL line isn't low after high phase");
	               end
	               
	               #(third*10);
	               //Transition to next bit
	           end
	           
	           /*Master is sending out ack or nack bits*/
	           else begin
	               sda_reg = 'z;
	               
	               #10;
	               
	               /*Master should have sent out nack bit*/
	               if(k == count-1) begin
	                   assert(SDA == '1) begin
	                   end else begin $display("Master hasn't sent out nack bit");
	                   end
	               end
	               
	               /*Master sends out ack bit*/
	               else begin
	                   assert(SDA == '0) begin
	                   end else begin $display("Master hasn't sent out ack bit");
	                   end
	               end 
	               
	               //In both cases SCL is low
	               assert(scl == '0) begin
	               end else begin $display("SCL should be low as master sends out ack/nack bit");
	               end
	               
	               #((third-1)*10);
	               
	               //Read 2 state
	               assert(SDA == (k == count - 1)) begin
	               end else begin 
	               $display("Slave has changed SDA control during SCL high phase");
	               end
	               
	               assert(scl == '1) begin
	               end else begin $display("SCL line isn't high");
	               end
	               
	               #(third*10);
	               //Read 3 state
	               assert(SDA == (k == count - 1)) begin
	               end else begin 
	               $display("Slave has changed SDA control during SCL low phase");
	               end
	               
	               assert(scl == '0) begin
	               end else begin $display("SCL line isn't low after high phase");
	               end
	               
	               #(third*10);
	               //Transition to next byte or to stop state
	           end  
	       end
	       k = k + 1;
	   end
	endtask
	
	logic[1:0][7:0] random_rx_byte;
	
	//STIMULUS BLOCK  
	initial begin
	   clk = '0;
	   
	    while($time < 2000000000) begin
	      sda_reg = 'z; //SDA has open drain structure with pullup resistors
		  /*Initialize i2cmaster*/
		  reset = '1;
		
		  #10;
		
		  /*Randomize inputs */
		  reset = '0;
		  randomized_inputs(valid_instr, full_i2cbuffer, wr_data, mode, reg_address);
		  
		  /*If appropriate signals aren't received*/
		  if(full_i2cbuffer || valid_instr[0] == '0) begin
		      
		      #2;
		      if (full_i2cbuffer) begin
		          assert(master_free == '0) begin
		          end else begin
		          $display("Master free for new transaction even when queue is full");
		          end
		      end
		      
		      #8;
		      continue;
		  end
		  
		  /*System in idle state.*/
		  #10;
		  /*System is in start 1 state. All future state transitions
		  take place after a third of an SCL clock period*/
		  
		  assert(controller.address_reg == reg_address) begin
		  end else begin $display("Register address not stored"); end
		  
		  assert(controller.valid_reg == valid_instr) begin
		  end else begin $display("Valid signals not stored"); end
		  
		  assert(controller.data_reg == wr_data) begin
		  end else begin $display("Data to write not stored"); end
		  
		  assert(controller.mode_reg == mode) begin
		  end else begin $display("Operation info not stored"); end
		  
		  assert(controller.hold_sda == 1'b1) begin
		  end else begin $display("SDA not held by master to initiate communication");
		  end
		  
		  assert(scl == '1) begin
		  end else begin $display("SCL line not held high by master before signalling start");
		  end
		  
		  
		  assert(scl == '1) begin
		  end else begin $display("SCL line not high when SDA is pulled low to signal start");
		  end
		  
		  assert(SDA == '0) begin
		  end else begin $display("SDA not pulled low to signal start");
		  end
		  $display($time);
		  
		  /*Transistion to start 2 state*/
		  #((third)*10); 
		  
		  assert(scl == '0) begin
		  end else begin $display("SCL not pulled low to signal start condition");
		  end
		  
		  assert(SDA == '0) begin
		  end else begin $display("SDA not pulled low to signal start condition");
		  end
		  
		  /*Transition to address 1 state*/
		  #((third)*10);
		  
		  write_vector = {serialbusaddr, 2'b0};
		  
		  //For transmitting serial bus address byte.
		  write_phase_check(write_vector,6);
		  
		  /*Transition into address 4 state*/
		  write_vector = {reg_address,1'b0};
		  write_phase_check(write_vector,5);
		  
		  /*Transition into write/read state*/
		  if(mode[2] || mode[3]) begin
		      /*If sending out 2 bytes of data,
		      start with most significant byte*/
		      if(mode[3]) begin
		          write_vector = {wr_data[15:8],1'b0};
		          write_phase_check(write_vector,4);
		          
		          /*Send out least significant byte*/
		          write_vector = {wr_data[7:0],1'b0};
		          write_phase_check(write_vector,3);
		      end
		      
		      
		      /*Otherwise if sending out 1 byte*/
		      else begin
		          write_vector = {wr_data[7:0],1'b0};
		          write_phase_check(write_vector,4);
		          /*Transition into stop state*/
		      end
		      
		      /*Or transition into stop state*/    
		  end
		  
		  else if(mode[0] || mode[1]) begin
		      read_phase_check(mode,random_rx_byte);
		      
		      /*Check to see if we received the correct data
		      for a 2 - byte read*/
		      if(mode[1]) begin
		          assert(controller.received_data == {random_rx_byte[1],random_rx_byte[0]}) 
		          begin end else 
		          begin 
		          $display("2 byte read data not registered appropriately");
		          end
		      end
		      
		      /*Check to see if correct byte ws received*/
		      else begin
		          assert(controller.received_data[7:0] == {random_rx_byte[1]}) 
		          begin end else 
		          begin 
		          $display("Single byte read data not registered appropriately");
		          end
		      end
		      
		      
		  end
		  
		  //Transitioned into stop state
		  assert(SDA == '0) begin end else begin 
		  $display("SDA hasn't transitioned to 0 to prepare to signal stop state");
		  end
		  
		  assert(scl == '0) begin end else begin
		  $display("scl not low when SDA transition to 0 to prepare to signal stop");
		  end
		  
		  #((third)*10);
		  //Stop State 2
		  assert(SDA == '0) begin end else begin
		  $display("SDA should be low during SCl high phase in stop state 2");
		  end
		  
		  assert(scl == '1) begin end else begin
		  $display("scl should be high during stop state 2");
		  end
		  
		  #(third*10);
		  //Stop State 3
		  assert(SDA == '1) begin end else begin
		  $display("SDA should have transitioned to high with scl high to signal stop");
		  end
		  
		  assert(scl == '1) begin end else begin
		  $display("scl should be high to during stop state 3");
		  end
		  
		  #((third-1)*10);
		  assert(i2c_data_rdy == '1) begin end else begin
		  $display("Controller hasn't signalled communication completion");
		  end
		  
		  #20;
		  //Wait for buffer to be written
		  #10;
		  //Transition to idle state at the end of the loop
	   end
	end
endmodule
	
	
