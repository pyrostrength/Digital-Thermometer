/*I2C master controller for the temperature sensor.

To read data from temperature sensor, communication operates
in the following format:
For 1-byte read:
Start -> Serial Bus Address Byte + Read -> Ack(from slave) -> Register Address
-> Ack(slave) -> Repeat Start -> Serial Bus Address + Read -> Ack(from slave) ->
Data Byte -> Nack(from Master) -> Stop

For 2-byte reads:
Start -> Serial Bus Address Byte + Read -> Ack(from slave) -> Register Address 
-> Ack(slave) -> Repeat Start -> Serial Bus Address + Read -> Ack(from slave) ->
Data Byte 1 -> Ack(from Master) -> Data Byte 2 -> Nack(from Master) -> Stop

For 1 byte writes:
Start -> Serial Bus Address Byte + Read -> Ack(from slave) -> Register Address 
-> Ack(slave) -> Data Byte 1 -> Ack(from slave) -> Stop

For 2 byte writes:
Start -> Serial Bus Address Byte + Read -> Ack(from slave) -> Register Address ->
Ack(slave) -> Data Byte 1 -> Ack(from slave) -> Data Byte 2 -> Ack(from slave)
-> Stop

All operations with ADT7420 are initiated in the form of read/writes.

Controller registers all instruction data necessary for operation and sends
it out to buffer in next pipeline stage when communication is complete.

In I2C communication data changes only during the low period of SCL clock. Therefore we sample
the data after SCL low phase but before the middle portion of the SCL high phase.
*/

module i2cmaster(input logic clk,reset,
                 /*If buffers on next pipeline stage are full,
                 we do not initiate communication*/
				 input logic full_i2cbuffer, 
				 input logic[15:0] wr_data,//Data to write to temp sensor registers
				 /*Operation to be performed. 1st 4 bits
				 are {write_2byte, write_1byte,read_2byte,read_1byte}*/
				 input logic[7:0] mode,
				 input logic[1:0] valid_instr,//signal to initiate I2C communication
				 input logic[6:0] serialbusaddr, //serial bus address for temp sensor
				 input logic[7:0] reg_address, //address of temperature sensor register
				 input logic[9:0] dvsr, //number of cycles of system clock per I2C clock cycle
				 output logic[15:0] received_data, //Data received from reading SDA line
				 output logic master_free, //Indicates controller is ready to initiate communication
				 output logic[5:0] failure_signal,//Indicates read/write failure
				 output logic i2c_data_rdy,//Indicates completion of communication
				 
				 /*Info for completed instruction to be passed onto next pipeline
				 stage*/
				 output logic[1:0] i2c_valid_instr,
				 output logic[15:0] i2c_retrieved_data,
				 output logic[7:0] i2c_op_info,
				 output logic[7:0] i2c_instr_address,
				 
				 output tri scl, //SCL clock generated by master
				 inout tri sda); //Serial Data Line.
				     
				        
				 typedef enum { 
				    idle,start1,start2, address1,address2,address3,address4,address5,address6,
				    restart1,restart2,restart3,restart4,
				    read1,read2,read3,read4,read5,read6,
				    write1,write2,write3,write4,write5,write6,
				    stop1,stop2,stop3} state_type;
				 
				 state_type state, state_next;
				 logic sda_reg, sda_next;
				 logic scl_reg, scl_next;
				 logic[9:0] count, count_next; //Counter for I2C clock cycle
				 logic[4:0] bit_reg,bit_next; //Counts number of bits transmitted or received.
				 logic[9:0] qutr,half; //Numbers corresponding to quarter and half of SCL clock cycle
				     	
				 logic write;
				 logic hold_sda,read_phase;
			     logic[8:0] write_reg, write_next; //Holds data to be written on SDA
			     
			     /*Since reads requires resending the serial bus address,
			     we make the state machine code more concise by having control
			     signals that determine whether we transition to reading data from SDA
			     after sending the serial bus address or if we transition to sending
			     the register address*/
				 logic readbyte_next,readbyte_reg; 
				 logic[15:0] received_data_next;
				 
				 /*Control signals to indicate communication failure 
				 during each stage of I2C communication
				 when necessary ack/nack bit isn't received/sent*/
				 logic sba_send_fail, address_send_fail, write_byte1_fail, write_byte2_fail, read_byte1_fail, read_byte2_fail;
				 logic sba_send_fail_next, address_send_fail_next, write_byte1_fail_next, write_byte2_fail_next, read_byte1_fail_next, read_byte2_fail_next;
				  
				 /*Register to hold data for necessary for communication*/
				 logic[7:0] mode_next,mode_reg;
				 logic[15:0] data_next,data_reg;
				 logic[7:0] address_next,address_reg;
				 logic[2:0] valid_next,valid_reg;
				 
				    	
				 assign failure_signal = {sba_send_fail, address_send_fail, write_byte1_fail, write_byte2_fail, read_byte1_fail, read_byte2_fail};
				 assign qutr = dvsr / 4;
				 assign half = dvsr /2;
				  	
				 always_ff @(posedge clk,posedge reset) begin
				    if(reset) begin
				        state <= idle;
				        sda_reg <= '1;
				     	scl_reg <= '1;
				     	bit_reg <= '0;
				     	count <= '0;
				     	received_data <= '0;
				     	write_reg <= '0;
				     	readbyte_reg <= '0; 
				     			
				     			
				     	sba_send_fail <= '0; 
				     	address_send_fail <= '0;
				     	write_byte1_fail <= '0;
				     	write_byte2_fail <= '0;
				     	read_byte1_fail <= '0;
				     	read_byte2_fail <= '0;
				     	
				     	i2c_valid_instr <= '0;
				     	i2c_retrieved_data <= '0;
				     	i2c_op_info <= '0;
				     	i2c_instr_address <= '0;
				     	
				     end
				     		
				     else begin
				     	received_data <= received_data_next;
				     	readbyte_reg <= readbyte_next;
				     	sda_reg <= sda_next;
				     	count <= count_next;
				     	scl_reg <= scl_next;
				     	state <= state_next;
				     	bit_reg <= bit_next;
				     	write_reg <= write_next;
				     			
				     	sba_send_fail <= sba_send_fail_next; 
				     	address_send_fail <= address_send_fail_next;
				     	write_byte1_fail <= write_byte1_fail_next;
				     	write_byte2_fail <= write_byte2_fail_next;
				     	read_byte1_fail <= read_byte1_fail_next;
				     	read_byte2_fail <= read_byte2_fail_next;
				     	
				     	valid_reg <= valid_next;
				     	data_reg <= data_next;
				     	mode_reg <= mode_next;
				     	address_reg <= address_next;
				     end
				 end
				 
				 /*SCL and SDA have open-drain structure.When not driven
				 the lines are pulled high.*/ 					   					
			     assign scl = (scl_reg) ? 1'bz: 1'b0;
					
			     /*If slave is driving sda line then output on master is in
			     high impedance state and SDA value depends on what
			     slave drives it to. If master is holding the SDA line and
			     requires to write 1 to it, then if output is high impedance
			     state then SDA line is pulled high*/	
				 assign sda = (read_phase || (hold_sda && sda_reg))? 1'bz : 1'b0; 
				 
				 /*During writes,Master only writes 8 bits to temperature sensor 
				 b4 receiving ack/nack bit. If Master is reading from temp sensor
				 then it only writes the ack/nack bit*/	
				 assign write = (hold_sda && (bit_reg < 8)) || (read_phase && (bit_reg == 8));
				 
				 assign i2c_valid_instr = valid_reg;
				 
				 assign i2c_retrieved_data = data_reg;
				 
				 assign i2c_op_info = mode_reg;
				 
				 assign i2c_instr_address = address_reg;
				 			
				 //State machine logic
				 always_comb begin
				    i2c_data_rdy = 1'b0;
				    state_next = state;
				    bit_next= bit_reg;
				    scl_next = 1'b1;
				    count_next = count + 1;
				    sda_next = write_reg[8];
				    hold_sda = 1'b0;
				    read_phase = 1'b0;
				    master_free = 1'b0;
				    write_next = write_reg; 
				    readbyte_next = readbyte_reg;
				    received_data_next = received_data;
				     		
				    //Failure signals need to be registered, otherwise they are lost
				    sba_send_fail_next = sba_send_fail; 
				    address_send_fail_next = address_send_fail;
				    write_byte1_fail_next = write_byte1_fail;
				    write_byte2_fail_next = write_byte2_fail;
				    read_byte1_fail_next = read_byte1_fail;
				    read_byte2_fail_next = read_byte2_fail;
				     
				    mode_next = mode_reg;
				    valid_next = valid_reg;
				    data_next = data_reg;
				    address_next = address_reg;
				    
				     		
				    case(state)
				        idle: begin
				     	  sda_next = 1'b1;
				     	  /*I2C controller cannot initiate communication
				     	  if buffers in next pipeline is full. So we
				     	  propagate the stall to prior stage in the pipeline
				     	  to prevent clearing of instruction from buffer*/
				     	  master_free = (!full_i2cbuffer);
				     	  
				     	  /*Communication can be initiated only if a valid instruction is
				     	  requesting communication and buffers on next stage of pipeline aren't
				     	  full.
				     	  Valid_instr[0] is high if an instruction made a request or under
				     	  default mode of operation*/
				     	  if(valid_instr[0] & full_i2cbuffer) begin 
				     	      state_next = start1;
				     		  sda_next = 1'b0;
				     		  count_next = '0;
				     		  /*We write the serial bus address to temp sensor
				     		  thus read segment of write_next == 1'b0 */
				     		  write_next = {serialbusaddr, 2'b0};
				     		  
				     		  //Store instruction data
				     		  mode_next = mode;
				     		  valid_next = valid_instr;
				     		  data_next = wr_data;
				     		  address_next = reg_address;
				     	  end
				        end
				     			
				     	start1: begin
				     	  hold_sda = 1'b1; //Hold sda and drive it low
				     	  sda_next = 1'b0;
				     	  /*Keep SCL high and drive SDA low to signal start
				     	  condition*/ 
				     	  scl_next = 1'b1; 
				     	  if(count == qutr - 1) begin
				     	      state_next = start2; 
				     		  count_next = '0;
				     		  scl_next = '0; 
				     	  end
				     	end
				     			
				     	start2:begin
				     	  hold_sda = 1'b1;
				     	  sda_next = '0; //Hold SCL and SDA low for quarter SCL clock cycle
				     	  scl_next = '0;
				     	  if(count == qutr - 1) begin
				     	      state_next = address1;
				     		  count_next = '0;
				     	  end
				     	end
				     			
				     	/*Write serial bus address byte identifying I2C temp sensor to SDA*/
				     	address1:begin
				     	  scl_next = 1'b0; 
				     	  hold_sda = 1'b1;
				     	  if(count == qutr - 1) begin
				     		  state_next = address2;
				     		  count_next = '0;
				     		  scl_next = 1'b1;  
				     	  end
				     	end
				     			
				     	/*Data has been read off SDA line at SCL positive clock edge*/
				     	address2:begin
				     	  hold_sda = 1'b1; 
				     	  scl_next = 1'b1;
				     	  if(count == qutr - 1) begin
				     	      received_data_next = (bit_reg != 8) ? {received_data[15:1], sda} : received_data;
				     	      sba_send_fail_next  = (bit_reg == 8 && sda != 0) ? 1'b1 : sba_send_fail;
				     	  end
				     	  if(count == half - 1) begin
				     	      scl_next = 1'b0;
				     		  state_next = address3;
				     		  count_next = '0;
				     	  end
				     	end
				     			
				     	address3: begin
				     	  hold_sda = 1'b1;
				     	  scl_next = 1'b0; //Hold scl low
				     	  if(count == qutr - 1) begin 
				     	      count_next = '0;
				     		  if(bit_reg == 8) begin //Data byte + ack/nack bit
				     		     bit_next = 1'b0;  //Reset bit counter
				     		     /*Proceed to reading off data byte after writing serial bus address byte 
				     		     or proceed with writing register address*/
				     			 state_next = (readbyte_reg) ? read1 : address4; 
				     			 write_next = (readbyte_reg) ? {9{mode_reg[0]}} : {address_reg,1'b0};
				     			 readbyte_next = '0;
				     		  end
				     					
				     		  //Some address bits haven't been transmitted 
				     		  else  begin 
				     		     state_next = address1; 
				     			 bit_next = bit_reg + 1'b1;
				     			 write_next = {write_reg[7:0], 1'b0};
				     		  end
				     	  end
				     	end
				     			
				     	/*Write register address to SDA*/
				     	address4:begin
				     	  scl_next = 1'b0; 
				     	  hold_sda = 1'b1;
				     	  if(count == qutr - 1) begin
				     		  state_next = address5;
				     		  count_next = '0;
				     		  scl_next = 1'b1;
				     	  end
				     	end
				     			
				     	address5:begin
				     	  hold_sda = 1'b1; 
				     	  scl_next = 1'b1; 
				     	  if(count == qutr - 1) begin
				     	      received_data_next = (bit_reg != 8) ? {received_data[15:1], sda} : received_data;
				     	      address_send_fail_next  = (bit_reg == 8 && sda != 0) ? 1'b1 : address_send_fail;
				     	  end
				     	  if(count == half - 1) begin
				     	      scl_next = 1'b0;
				     		  state_next = address6;
				     		  count_next = '0;
				     	  end
				     	end
				     			
				        /*From this state,transition to either reading or writing from/to the SDA*/
				     	address6: begin
				     	  hold_sda = 1'b1;
				     	  scl_next = 1'b0; 
				     	  if(count == qutr - 1) begin 
				     	      count_next = '0;
				     		  if(bit_reg == 8) begin
				     		     bit_next = 1'b0;
				     			 if(mode_reg[0] || mode_reg[1]) begin
				     			    state_next = restart1;
				     				write_next = 9'b0;
				     			 end
				     			 
				     			 else if(mode_reg[2] || mode_reg[3])  begin
				     			    state_next = write1;
				     			    /*If we need only write 1 byte, otherwise...*/
				     			    /*In 2 byte write M.S.Byte sent out first*/
				     				write_next = (mode_reg[2]) ? {data_reg[7:0], 1'b0} : {data_reg[15:8], 1'b0};
				     			 end
				     						
				     			 else begin
				     			    state_next = stop1;
				     			 end
				     		  end
				     					
				     		  //Some address bits haven't been transmitted 
				     		  else  begin 
				     		     state_next = address4; 
				     			 write_next = {write_reg[7:0], 1'b0};
				     			 bit_next = bit_reg + 1'b1;
				     		  end
				     	   end
				        end
				     			
				     	/*Writing to I2C temperature sensor*/
				     	write1: begin
				     	  scl_next = '0;
				     	  hold_sda = 1'b1;
				     	  if(count == qutr - 1) begin
				     		  state_next = write2;
				     		  count_next = '0;
				     		  scl_next = 1'b1;
				     	  end
				     	end
				     	
				     			
				     	write2: begin
				     	  hold_sda = 1'b1;
				     	  scl_next = 1'b1;
				     	  if(count == qutr - 1) begin
				     	      received_data_next = (bit_reg != 8) ? {received_data[15:1], sda} : received_data;
				     	      write_byte1_fail_next  = (bit_reg == 8 && sda != 0) ? 1'b1 : write_byte1_fail;
				     	  end
				     	  if(count == half-1) begin
				     	      scl_next = 1'b0;
				     		  state_next = write3;
				     		  count_next = '0;
				     	  end
				     	end
				     			
				     	write3:begin
				     	  hold_sda = 1'b1;
				     	  scl_next = 1'b0; //Hold scl low
				     	  if(count == qutr-1) begin 
				     	      count_next = '0;
				     		  if(bit_reg == 8) begin //Data byte + ack/nack bit
				     		     bit_next = 1'b0;
				     			 /*If we're writing 2 bytes of data*/
				     			 if(mode_reg[3]) begin
				     			    state_next = write4;
				     				write_next = {data_reg[7:0],1'b0};
				     			 end
				     						
				     			 //Finished writing the necessary data
				     			 else begin
				     			    state_next = stop1;
				     			 end
				     		  end
				     		  //Write is incomplete.
				     		  else  begin
				     		     write_next = {write_reg[7:0], 1'b0};
				     			 state_next = write1; 
				     			 bit_next = bit_reg + 1'b1;
				     		  end
				     	  end
				     	end
				     			
				     	/*Writing 2nd byte*/
				     	write4: begin
				     	  scl_next = '0;
				     	  hold_sda = 1'b1;
				     	  if(count == qutr-1) begin
				     		  state_next = write5;
				     		  count_next = '0;
				     		  scl_next = 1'b1;
				     	  end
				     	end
				     			
				     	write5: begin
				     	  hold_sda = 1'b1;
				     	  scl_next = 1'b1; //Hold scl high.
				     	  if(count == qutr - 1) begin
				     	      received_data_next = (bit_reg != 8) ? {received_data[15:1], sda} : received_data;
				     	      write_byte2_fail_next  = (bit_reg == 8 && sda != 0) ? 1'b1 : write_byte2_fail;
				     	  end
				     	  if(count == half-1) begin
				     	      scl_next = 1'b0;
				     		  state_next = write6;
				     		  count_next = '0;
				     	  end
				     	end
				     			
				     	write6:begin
				     	  hold_sda = 1'b1;
				     	  scl_next = 1'b0; //Hold scl low
				     	  if(count == qutr-1) begin 
				     	      count_next = '0;
				     		  if(bit_reg == 8) begin //Data byte + ack/nack bit
				     		     bit_next = 1'b0; 
				     		     state_next = stop1;
				     		  end
				     					
				     		  //Write is incomplete.
				     		  else  begin
				     		     write_next = {write_reg[7:0],1'b0};
				     			 state_next = write4; 
				     			 bit_next = bit_reg + 1;
				     		  end
				     	  end
				     	end
				     				
				     			
				     	/*Initiate repeat start by pulling sda high*/
				        restart1:begin
				     	  scl_next = 1'b0;
				     	  sda_next = 1'b1;
				     	  hold_sda = '1;
				     	  if(count == qutr - 1) begin
				     	      scl_next = 1'b1;
				     		  count_next = '0;
				     		  state_next = restart2;
				     	  end
				     	end
				     			
				     	//SCL high. We initiate SDA transition during the midpoint of SCL's high phase.
				        restart2:begin
				          hold_sda = '1;
				     	  scl_next = 1'b1;
				     	  sda_next =  1'b1;
				     	  if(count == qutr - 1) begin
				     	      state_next = restart3;
				     		  count_next = '0;
				     		  sda_next = '0; 
				     	  end
				     	end
				     			
				     	restart3:begin
				     	  hold_sda = '1;
				     	  scl_next = 1'b1;
				     	  sda_next = 1'b0;
				     	  if(count == qutr - 1) begin
				     	      state_next = restart4;
				     		  scl_next = 1'b0;
				     		  count_next = '0;
				     	  end
				     	end

				     	restart4:begin
				     	  scl_next = 1'b0;
				     	  sda_next = 1'b0;
				     	  if(count == qutr - 1) begin
				     	      state_next = address1;
				     		  scl_next = 1'b0;
				     		  count_next = '0;
				     		  readbyte_next = 1'b1;
				     		  /*The 1'b1 is necessary since we need to indicate
				     		  to temp sensor that we're reading from it*/
				     		  write_next = {serialbusaddr , 1'b1, 1'b0};
				     	  end
				     	end
				     			
				     	read1: begin
				     	  scl_next = '0;
				     	  read_phase = 1'b1;
				     	  if(count == qutr - 1) begin
				     		  state_next = read2;
				     		  count_next = '0;
				     		  scl_next = 1'b1;
				     	  end
				     	end
				     			
				     	read2: begin
				            read_phase = 1'b1;
				     		scl_next = 1'b1; //Hold scl high.
				     		if(count == qutr - 1) begin
				     	      received_data_next = (bit_reg != 8) ? {received_data[15:1], sda} : received_data;
				     	      read_byte1_fail_next  = (bit_reg == 8 && sda != 0) ? 1'b1 : read_byte1_fail;
				     	    end
				     		
				     		if(count == half - 1) begin
				     		 scl_next = 1'b0;
				     		 state_next = read3;
				     		 count_next = '0;
				     		end
				     	end
				     			
				     			
				     	read3:begin
				     	  read_phase = 1'b1;
				     	  scl_next = 1'b0; //Hold scl low
				     	  if(count == qutr - 1) begin 
				     	      count_next = '0;
				     		  if(bit_reg == 8) begin //Data byte + ack/nack bit
				     		     bit_next = 1'b0;
				     		     /*If reading 2 bytes*/ 
				     			 if(mode_reg[1]) begin
				     			    state_next = read4;
				     			    /*Master must send a nack bit
				     			    to acknowledge receiving final bit.Nack bit is 1*/
				     				write_next = {9{mode_reg[1]}};
				     			 end
				     						
				     			 else begin
				     			    state_next = stop1;
				     			 end	
				     	      end
				     						
				     	      //Read is incomplete. Perform shifing on write data to get to the ack/nack bit
				     	      else  begin
				     	         state_next = read1; 
				     		     bit_next = bit_reg + 1'b1;
				     		     write_next = {write_reg[7:0],1'b0};
				     	      end
				           end
				        end
				     			
				     	read4: begin
				     	  scl_next = '0;
				     	  read_phase = 1'b1;
				     	  if(count == qutr - 1) begin
				     		  state_next = read5;
				     		  count_next = '0;
				     		  scl_next = 1'b1;
				     	  end
				     	end
				     	
				     	read5: begin
				     	  read_phase = 1'b1; //Data has been shifted in at clock edge of state transition from address1 to address2
				     	  scl_next = 1'b1; //Hold scl high.
				     	  
				     	  if(count == qutr - 1) begin
				     	      received_data_next = (bit_reg != 8) ? {received_data[15:1], sda} : received_data;
				     	      read_byte2_fail_next  = (bit_reg == 8 && sda != 1) ? 1'b1 : read_byte2_fail;
				     	  end
				     	  
				     	  if(count == half - 1) begin
				     	      scl_next = 1'b0;
				     		  state_next = read6;
				     		  count_next = '0;
				     	  end
				     	end
				     			
				     			
				     	read6:begin
				     	  read_phase = 1'b1;
				     	  scl_next = 1'b0; //Hold scl low
				     	  if(count == qutr - 1) begin 
				     	      count_next = '0;
				     		  if(bit_reg == 8) begin //Data byte + ack/nack bit
				     		     bit_next = 1'b0; 
				     			 state_next = stop1;
				     			 //SDA must be pulled low in preparation of pulling
				     			 //it high when SCL is high to signal stop 
				     			 sda_next = '0; 
				     		  end
				     					
				     		  else  begin
				     		     state_next = read4; 
				     			 bit_next = bit_reg + 1'b1;
				     			 write_next = {write_reg[7:0],1'b0};
				     		  end
				     	  end
				     	end
				     			
		
				     	/*SDA is pulled low*/
				     	stop1:begin
				     	  scl_next = '0;
				     	  sda_next = '0;
				     	  hold_sda = 1'b1;
				     	  if(count == qutr - 1) begin
				     	      state_next = stop2;
				     		  count_next = '0;
				     		  scl_next = 1'b1;
				     	  end
				     	end
				     			
				     	stop2:begin
				     	  scl_next = 1'b1;
				     	  sda_next = 1'b0;
				     	  hold_sda = 1'b1;
				     	  if(count == qutr - 1) begin
				     	      state_next = stop3;
				     		  count_next = '0;
				     		  sda_next = '1;
				     	  end
				     	end
				     			
				     	/*SDA to high and hold for a quarter cycle before transitioning to idle state*/
				     	stop3:begin
				     	  hold_sda = 1'b1;
				     	  scl_next = 1'b1;
				     	  sda_next = 1'b1;
				     	  if(count == qutr -1) begin
				     	      state_next = idle;
				     		  count_next = '0;
				     		  i2c_data_rdy = 1'b1;
				     	  end
				     	end
							
				   endcase
		         end			
endmodule
				     				
				     					
				     				
				     					
				     				
				     				
				     			
				     				
				     				
				     				
				     				
				     					
				     					
				     				
				     				
				     					
				     					
				     					
				     			
				     			
				     		
				     		
				     	
				     	
				     	
				     		
				     		
				     	
				     	
				     	
					
				     
				  
