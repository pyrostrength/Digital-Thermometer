/*I2c controller works for reading and writing bytes to i2c temp sensor*/

module i2cmaster_test ;

	logic clk,reset;
	logic[15:0] wr_data;
	logic[2:0] mode; //read 1/2 bytes, write 1/2 bytes, general call and reset.
	logic initiate; //signal from processor/driver to initiate I2C transaction
	logic[6:0] serialbusaddr;//serial bus address for the temp sensor 
	logic[7:0] addrpointer; //address pointer byte for specific register to access
	logic[9:0] dvsr; //number of cycles of "clk" per I2C clock cycle
	logic[15:0] received_data;//Receiving shift register that stores reads off of the sda line.
	logic ready; //indicates master is available for an I2C transaction
	tri scl; //SCL clock generated by master
	tri sda;//SDA line
	
	logic SDA; //Secondary sda line for implementing open drain structure of SDA line in I2C comms
	
	i2cmaster controller(.clk(clk),
						 .sda(sda),
						 .scl(scl),
						 .ready(ready),
						 .received_data(received_data),
						 .dvsr(dvsr),
						 .addrpointer(addrpointer),
						 .serialbusaddr(serialbusaddr),
						 .initiate(initiate),
						 .wr_data(wr_data),
						 .mode(mode),
						 .reset(reset));
	
	assign SDA = (sda === 1'bz)? 1'b1:sda;
	
	`timescale 1ns/1ps
	
	always begin
		#5 clk = ~clk;
	end
	
	initial begin
		/*Initialize i2cmaster by reset*/
		clk = '0;
		reset = 1'b1;
		
		#10;
		/*Initiate writing of 1 byte*/
		reset = '0;
		serialbusaddr = 7'b1011101;
		addrpointer = 8'b00000010;
		wr_data = 8'b01011101;
		mode = 3'b010;
		dvsr = 10'b00000_01000; //Nothing happens. No initiate signal given.
		
		#10
		initiate = 1'b1; //Now we initiate the writing of 1 byte.
		
		#50 //We need to transition completely out of idle state so that...
		initiate = 1'b0;
		
		wait(ready == 1'b1); //when we complete writing a byte we test for writing 2 bytes:)
		initiate = 1'b1;
		mode = 3'b011; //Writing 2 bytes
		wr_data = 16'b00101011_01101100;
		
		#50
		initiate = 1'b0;
		
		wait(ready == 1'b1); //We shall now test for reading 1 byte or 2 bytes. Then we design UART CORE :);
		initiate = 1'b1;
		mode = 3'b000; //Test for reading 1 byte
		
		#50
		wait(ready == 1'b1);
		mode = 3'b001; //Test for reading 2 byte
		
	end
endmodule
	
	
