module i2c_uart_arbiter_tb;
endmodule
