//Minimum I2C clock rate is 8 system clock cycles per I2C clock cycle.
//Avoiding prior setup limits the overall clock speed.
//Clock speed relatively slow - speed at 150MHz.

module i2cmaster (input logic clk,reset,
				     input logic[15:0] wr_data,
				     input logic[2:0] mode, //read 1/2 bytes, write 1/2 bytes, general call and reset.
				     input logic initiate, //signal from processor/driver to initiate I2C transaction
				     input logic[6:0] serialbusaddr, //serial bus address for temp sensor
				     input logic[7:0] addrpointer, //address pointer byte for specific register to access
				     input logic[9:0] dvsr, //number of cycles of "clk" per I2C clock cycle
				     output logic[15:0] received_data, //Receiving shift register that stores reads off of the sda line.
				     output logic ready, //indicates master is available for an I2C transaction
				     output tri scl, //SCL clock generated by master
				     inout tri sda); //Serial Data Line.
				     
				        
				        typedef enum { 
				     	idle,start1,start2, address1,address2,address3,address4,address5,address6,
				     	restart1,restart2,restart3,restart4,
				     	read1,read2,read3,read4,read5,read6,
				     	write1,write2,write3,write4,write5,write6,
				     	stop1,stop2,stop3} state_type;
				     
				     
				     	state_type state, state_next;
				     	logic sda_reg, sda_next;
				    	logic scl_reg, scl_next;
				     	logic[9:0] count, count_next; //Counter for I2C clock cycle
				     	logic[4:0] bit_reg,bit_next; //Counting number of bits transmitted or received.
				     	logic[9:0] qutr,half; //count for dividing I2C/SCL clock cycle into 4 phases
				     	logic transmit_tick;
				     	
				     	logic write;
				     	logic hold_sda,read_phase;
					logic[8:0]write_reg, write_next;
					logic read_cmd, write_cmd,write2_cmd,read2_cmd;
					logic readbyte_next,readbyte_reg;
					logic[15:0] received_data_next;
				     	
				     	
				    	assign qutr = dvsr / 4;
				   	assign half = dvsr /2;
				   	
				   //Write, read and address states are identical in logic. Can condense them into one. Don't give up . Think. 
				   //Next state logic
				     always_ff @(posedge clk,posedge reset) begin
				     		if(reset) begin
				     			state <= idle;
				     			sda_reg <= '1;
				     			scl_reg <= '1;
				     			bit_reg <= '0;
				     			count <= '0;
				     			received_data <= '0;
				     			write_reg <= '0;
				     			readbyte_reg <= '0; 
				     			received_data <= '0;//Control signal simplifies state machine for reading a value. Need not add three more states
				     		end
				     		
				     		else begin
				     			received_data <= received_data_next;
				     			readbyte_reg <= readbyte_next;
				     			sda_reg <= sda_next;
				     			count <= count_next;
				     			scl_reg <= scl_next;
				     			state <= state_next;
				     			bit_reg <= bit_next;
				     			write_reg <= write_next;
				     		end
				     	end
				     					   					
					//assign scl = (scl_reg) ? 1'bz: 1'b0;
					
					assign scl = scl_reg;
					
					assign sda = (write)? sda_reg : 1'bz; 
					
					//assign sda = (!write || sda_reg) ? 1'bz : 1'b0;
					
					assign write = (hold_sda && (bit_reg < 8)) || (read_phase && (bit_reg == 8));
					
					always_comb begin
						read_cmd = 1'b0;
						write_cmd = 1'b0;
						read2_cmd = 1'b0;
						write2_cmd = 1'b0;
						case(mode)
							3'b000: begin
								read_cmd = 1'b1;
							end
							3'b001:begin
								read2_cmd = 1'b1;
							end
							3'b010:begin
								write_cmd = 1'b1;
							end
							3'b011:begin
								write2_cmd = 1'b1;
							end
						endcase
					end
								
				     	
				     	//State machine logic
				     	always_comb begin
				     		state_next = state;
				     		bit_next= bit_reg;
				     		scl_next = 1'b1;
				     		count_next = count + 1'b1;
				     		sda_next = write_reg[8];
				     		hold_sda = 1'b0;
				     		read_phase = 1'b0;
				     		ready = 1'b0;
				     		write_next = write_reg; 
				     		readbyte_next = readbyte_reg;
				     		received_data_next = received_data;
				     		
				     		case(state)
				     			idle: begin
				     				sda_next = 1'b1;
				     				ready = 1'b1;
				     				if(initiate) begin //We initiate a transaction.
				     					state_next = start1;
				     					sda_next = 1'b0;
				     					count_next = '0;
				     					write_next = {serialbusaddr, (write_cmd||write2_cmd), 1'b0};
				     				end
				     			end
				     			
				     			start1: begin
				     			    hold_sda = 1'b1; //Make and hold sda low.
				     				sda_next = 1'b0; 
				     				scl_next = 1'b1;
				     				if(count == qutr -1'b1) begin
				     					state_next = start2; 
				     					count_next = '0;
				     					scl_next = '0; //Make SCL low on next clock cycle/state transition
				     				end
				     			end
				     			
				     			start2:begin
				     			    hold_sda = 1'b1;
				     				sda_next = '0; //Hold SCL and SDA low for quarter SCL clock cycle
				     				scl_next = '0;
				     				if(count == qutr - 1'b1) begin
				     					state_next = address1;
				     					count_next = '0;
				     				end
				     			end
				     			
				     			/*Write serial bus address byte identifying I2C temp sensor to SDA*/
				     			address1:begin
				     				scl_next = 1'b0; 
				     				hold_sda = 1'b1;
				     				if(count == qutr-1'b1) begin
				     					state_next = address2;
				     					count_next = '0;
				     					scl_next = 1'b1;
				     					received_data_next ={received_data[15:1], sda};
				     				end
				     			end
				     			
				     			/*Data has been read off SDA line at SCL positive clock edge*/
				     			address2:begin
				     				hold_sda = 1'b1; 
				     				scl_next = 1'b1; 
				     				if(count == half-1'b1) begin
				     					scl_next = 1'b0;
				     					state_next = address3;
				     					count_next = '0;
				     				end
				     			end
				     			
				     			address3: begin
				     				hold_sda = 1'b1;
				     				scl_next = 1'b0; //Hold scl low
				     				if(count == qutr-1'b1) begin 
				     					count_next = '0;
				     					if(bit_reg == 8) begin //Data byte + ack/nack bit
				     						bit_next = 1'b0;  //Reset bit counter
				     						state_next = (readbyte_reg) ? read1 : address4; /*Proceed to reading off data byte after writing serial bus address byte or proceed with writing address pointer register byte*/
				     						write_next = (readbyte_reg) ? {9{read_cmd}} : {addrpointer,1'b0};
				     						//If write_cmd is 1, we write. If write_cmd is 0 then we read.
				     						readbyte_next = '0;
				     					end
				     					
				     					//Some address bits haven't been transmitted 
				     					else  begin 
				     						state_next = address1; 
				     						bit_next = bit_reg + 1'b1;
				     						write_next = {write_reg[7:0], 1'b0};
				     					end
				     				end
				     			end
				     			
				     			/*Write address pointer register byte to SDA*/
				     			address4:begin
				     				scl_next = 1'b0; 
				     				hold_sda = 1'b1;
				     				if(count == qutr-1'b1) begin
				     					state_next = address5;
				     					count_next = '0;
				     					scl_next = 1'b1;
				     					received_data_next ={ received_data[15:1], sda};
				     				end
				     			end
				     			
				     			address5:begin
				     				hold_sda = 1'b1; 
				     				scl_next = 1'b1; 
				     				if(count == half-1'b1) begin
				     					scl_next = 1'b0;
				     					state_next = address6;
				     					count_next = '0;
				     				end
				     			end
				     			
				     			/*From this state, transition to either reading or writing from/to the SDA*/
				     			address6: begin
				     				hold_sda = 1'b1;
				     				scl_next = 1'b0; 
				     				if(count == qutr-1'b1) begin 
				     					count_next = '0;
				     					if(bit_reg == 8) begin
				     						bit_next = 1'b0;
				     						if(read_cmd || read2_cmd) begin
				     							state_next = restart1;
				     							write_next = 9'b0;
				     						end
				     						
				     						else if(write_cmd || write2_cmd)  begin
				     							state_next = write1;
				     							write_next = (write_cmd) ? {wr_data[7:0], 1'b0} : {wr_data[15:8], 1'b0};
				     						end
				     						
				     						else begin
				     							state_next = stop1;
				     						end
				     						
				     					end
				     					
				     					//Some address bits haven't been transmitted 
				     					else  begin 
				     						state_next = address4; 
				     						write_next = {write_reg[7:0], 1'b0};
				     						bit_next = bit_reg + 1'b1;
				     					end
				     				end
				     			end
				     			
				     			/*Writing to I2C temperature sensor*/
				     			write1: begin
				     				scl_next = '0;
				     				hold_sda = 1'b1;
				     				if(count == qutr-1'b1) begin
				     					state_next = write2;
				     					count_next = '0;
				     					scl_next = 1'b1;
				     					received_data_next ={ received_data[15:1], sda};
				     				end
				     			end
				     			
				     			write2: begin
				     				hold_sda = 1'b1; //Data has been shifted in at clock edge of state transition from address1 to address2
				     				scl_next = 1'b1; //Hold scl high.
				     				if(count == half-1) begin
				     					scl_next = 1'b0;
				     					state_next = write3;
				     					count_next = '0;
				     				end
				     			end
				     			
				     			write3:begin
				     				hold_sda = 1'b1;
				     				scl_next = 1'b0; //Hold scl low
				     				if(count == qutr-1'b1) begin 
				     					count_next = '0;
				     					if(bit_reg == 8) begin //Data byte + ack/nack bit
				     						bit_next = 1'b0;
				     						/*If we're writing 2 bytes of data*/
				     						if(write2_cmd) begin
				     							state_next = write4;
				     							write_next = {wr_data[7:0],1'b0};//We shift out the lower byte in next clock cycle
				     						end
				     						
				     						//Finished writing the necessary data
				     						else begin
				     							state_next = stop1;
				     						end
				     					end
				     					
				     					//Write is incomplete.
				     					else  begin
				     						write_next = {write_reg[7:0], 1'b0};
				     						state_next = write1; 
				     						bit_next = bit_reg + 1'b1;
				     					end
				     				end
				     			end
				     			
				     			/*Writing 2nd byte*/
				     			write4: begin
				     				scl_next = '0;
				     				hold_sda = 1'b1;
				     				if(count == qutr-1'b1) begin
				     					state_next = write5;
				     					count_next = '0;
				     					scl_next = 1'b1;
				     					received_data_next ={ received_data[15:1], sda};
				     				end
				     			end
				     			
				     			write5: begin
				     				hold_sda = 1'b1;//Data has been shifted in at clock edge of state transition from address1 to address2
				     				scl_next = 1'b1; //Hold scl high.
				     				if(count == half-1) begin
				     					scl_next = 1'b0;
				     					state_next = write6;
				     					count_next = '0;
				     				end
				     			end
				     			
				     			write6:begin
				     				hold_sda = 1'b1;
				     				scl_next = 1'b0; //Hold scl low
				     				if(count == qutr-1'b1) begin 
				     					count_next = '0;
				     					if(bit_reg == 8) begin //Data byte + ack/nack bit
				     						bit_next = 1'b0; 
				     						state_next = stop1;
				     					end
				     					
				     					//Write is incomplete.
				     					else  begin
				     						write_next = {write_reg[7:0],1'b0};
				     						state_next = write4; 
				     						bit_next = bit_reg + 1'b1;
				     					end
				     				end
				     			end
				     				
				     			
				     			/*Initiate repeat start by pulling sda high*/
				     			restart1:begin
				     				scl_next = 1'b0;
				     				sda_next = 1'b1;
				     				if(count == qutr -1'b1) begin
				     					scl_next = 1'b1;
				     					count_next = '0;
				     					state_next = restart2;
				     				end
				     			end
				     			
				     			//SCL high. We initiate SDA transition during the midpoint of SCL's high phase.
				     			restart2:begin
				     				scl_next = 1'b1;
				     				sda_next =  1'b1;
				     				if(count==qutr-1'b1) begin
				     					state_next = restart3;
				     					count_next = '0;
				     				end
				     			end
				     			
				     			restart3:begin
				     				scl_next = 1'b1;
				     				sda_next = 1'b0;
				     				if(count == qutr -1'b1) begin
				     					state_next = restart4;
				     					scl_next = 1'b0;
				     					count_next = '0;
				     				end
				     			end
				     			
				     			restart4:begin
				     				scl_next = 1'b0;
				     				sda_next = 1'b0;
				     				if(count == qutr -1'b1) begin
				     					state_next = address1;
				     					scl_next = 1'b0;
				     					count_next = '0;
				     					readbyte_next = 1'b1;
				     					write_next = {serialbusaddr , 1'b0};
				     				end
				     			end
				     			
				     			read1: begin
				     				scl_next = '0;
				     				read_phase = 1'b1;
				     				if(count == qutr-1'b1) begin
				     					state_next = read2;
				     					count_next = '0;
				     					scl_next = 1'b1;
				     					received_data_next ={ received_data[15:1], sda};
				     				end
				     			end
				     			
				     			read2: begin
				     				read_phase = 1'b1;//Data has been shifted in at clock edge of state transition from address1 to address2
				     				scl_next = 1'b1; //Hold scl high.
				     				if(count == half-1'b1) begin
				     					scl_next = 1'b0;
				     					state_next = read3;
				     					count_next = '0;
				     				end
				     			end
				     			
				     			
				     			read3:begin
				     				read_phase = 1'b1;
				     				scl_next = 1'b0; //Hold scl low
				     				if(count == qutr-1'b1) begin 
				     					count_next = '0;
				     					if(bit_reg == 8) begin //Data byte + ack/nack bit
				     						bit_next = 1'b0; 
				     						if(read2_cmd) begin
				     							state_next = read4;
				     							write_next = {9{read2_cmd}};
				     						end
				     						
				     						else begin
				     							state_next = stop1;
				     						end	
				     					end
				     						
				     					//Read is incomplete. Perform shifing on write data to get to the ack/nack bit
				     					else  begin
				     						state_next = read1; 
				     						bit_next = bit_reg + 1'b1;
				     						write_next = {write_reg[7:0],1'b0};
				     					end
				     				end
				     			end
				     			
				     			read4: begin
				     				scl_next = '0;
				     				read_phase = 1'b1;
				     				if(count == qutr-1'b1) begin
				     					state_next = read5;
				     					count_next = '0;
				     					scl_next = 1'b1;
				     				end
				     			end
				     			
				     			read5: begin
				     				read_phase = 1'b1; //Data has been shifted in at clock edge of state transition from address1 to address2
				     				scl_next = 1'b1; //Hold scl high.
				     				if(count == half-1'b1) begin
				     					scl_next = 1'b0;
				     					state_next = read6;
				     					count_next = '0;
				     				end
				     			end
				     			
				     			
				     			read6:begin
				     				read_phase = 1'b1;
				     				scl_next = 1'b0; //Hold scl low
				     				
				     				if(count == qutr-1'b1) begin 
				     					count_next = '0;
				     					if(bit_reg == 8) begin //Data byte + ack/nack bit
				     						bit_next = 1'b0; 
				     						state_next = stop1;
				     					end
				     						
				     			
				     					else  begin
				     						state_next = read4; 
				     						bit_next = bit_reg + 1'b1;
				     						write_next = {write_reg[7:0],1'b0};
				     					end
				     				end
				     			end
				     			
		
				     			/*SDA is pulled low*/
				     			stop1:begin
				     				scl_next = '0;
				     				sda_next = '0;
				     				hold_sda = 1'b1;
				     				if(count == qutr - 1'b1) begin
				     					state_next = stop2;
				     					count_next = '0;
				     					scl_next = 1'b1;
				     				end
				     			end
				     			
				     			stop2:begin
				     				scl_next = 1'b1;
				     				sda_next = 1'b0;
				     				hold_sda = 1'b1;
				     				if(count == qutr -1'b1) begin
				     					state_next = stop3;
				     					count_next = '0;
				     				end
				     			end
				     			
				     			
				     			 /*SDA to high and hold for a quarter cycle before transitioning to idle state*/
				     			stop3:begin
				     				hold_sda = 1'b1;
				     				scl_next = 1'b1;
				     				sda_next = 1'b1;
				     				if(count == qutr -1'b1) begin
				     					state_next = idle;
				     					count_next = '0;
				     				end
				     			end
							
				     		endcase
				     	end
				
endmodule
				     				
				     					
				     				
				     					
				     				
				     				
				     			
				     				
				     				
				     				
				     				
				     					
				     					
				     				
				     				
				     					
				     					
				     					
				     			
				     			
				     		
				     		
				     	
				     	
				     	
				     		
				     		
				     	
				     	
				     	
					
				     
				  
